LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CLASS_32160462_MT IS


PORT(
	A, B : IN STD_LOGIC_VECTOR(1 downto 0);
	C : OUT STD_LOGIC_VECTOR(3 downto 0)
);
END CLASS_32160462_MT;

ARCHITECTURE MT_SYSTEM OF CLASS_32160462_MT IS

	COMPONENT CLASS_32160203_HA IS
	PORT(
	A,B:IN STD_LOGIC;
	S,C:OUT STD_LOGIC
	);
	END COMPONENT;
	
	SIGNAL REG_AND : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL REG_C : STD_LOGIC_VECTOR(3 downto 0);
	SIGNAL RES_SUM : STD_LOGIC;
	
BEGIN

	REG_AND(0) <= A(0) and B(0);
	REG_AND(1) <= A(0) and B(1);
	REG_AND(2) <= A(1) and B(0);
	REG_AND(3) <= A(1) and B(1);
	
	U1_HA : CLASS_32160203_HA
	PORT MAP(
		A=>REG_AND(1),
		B=>REG_AND(2),
		S=>REG_C(1),
		C=>RES_SUM
	);
	
	U2_HA : CLASS_32160203_HA
	PORT MAP(
		A=>RES_SUM,
		B=>REG_AND(3),
		S=>REG_C(2),
		C=>REG_C(3)
	);
	
	REG_C(0) <= REG_AND(0);
	C <= REG_C;
END MT_SYSTEM;