ENTITY half_adder IS
PORT(
	A,B:IN BIT;
	S,C:OUT BIT
);
END half_adder;

ARCHITECTURE ADDER OF half_adder IS
BEGIN

PROCESS(A,B)
BEGIN
	IF A=B THEN
		S<='0';
	ELSE
		S<='1';
	END IF;
END PROCESS;

PROCESS(A,B)
BEGIN
	IF A = '1' AND B = '1' THEN
		C<='1';
	ELSE
		C<='0';
	END IF;
END PROCESS;

END ADDER;
